version https://git-lfs.github.com/spec/v1
oid sha256:b266a9dd5394d8efa0e1eea8c4e631f8bfe9ee1004598a7f4545d486d8c00f73
size 8192
