version https://git-lfs.github.com/spec/v1
oid sha256:e96dce0db0d9a774ba9e3411e3bb4bf1be64793c866f21be36264a50c48ac926
size 3146240
